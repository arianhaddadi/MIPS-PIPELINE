module InstructionMem(input [31:0] address, output [31:0] instruction);
  reg [31:0] instructions [16383:0];
  integer i;
  initial begin
    for (i = 0 ; i <= 16383 ; i = i + 1) instructions[i] = {6'b000000, 26'b0};
		  instructions[0] = 32'b10001100000000010000001111101000;// lw r1,r0,1000
	    instructions[1] = 32'b00000000011000010001000000101010;// slt r2,r3,r1
	    instructions[2] = 32'b00000000000000000000000000000000;// nop
	    instructions[3] = 32'b00010000000000100000000000000001;// beq r2,r0,1
	    instructions[4] = 32'b00000000000000010001100000100000;// add r3,r1,r0
	    
	    instructions[5] = 32'b10001100000000010000001111101001;// lw r1,r0,1001
	    instructions[6] = 32'b00000000011000010001000000101010;// slt r2,r3,r1
	    instructions[7] = 32'b00000000000000000000000000000000;// nop
	    instructions[8] = 32'b00010000000000100000000000000001;// beq r2,r0,1
	    instructions[9] = 32'b00000000000000010001100000100000;// add r3,r1,r0
	    
	    instructions[10] = 32'b10001100000000010000001111101010;// lw r1,r0,1002
	    instructions[11] = 32'b00000000011000010001000000101010;// slt r2,r3,r1
	    instructions[12] = 32'b00000000000000000000000000000000;// nop
	    instructions[13] = 32'b00010000000000100000000000000001;// beq r2,r0,1
	    instructions[14] = 32'b00000000000000010001100000100000;// add r3,r1,r0
	    
	    instructions[15] = 32'b10001100000000010000001111101011;// lw r1,r0,1003
	    instructions[16] = 32'b00000000011000010001000000101010;// slt r2,r3,r1
	    instructions[17] = 32'b00000000000000000000000000000000;// nop
	    instructions[18] = 32'b00010000000000100000000000000001;// beq r2,r0,1
	    instructions[19] = 32'b00000000000000010001100000100000;// add r3,r1,r0
	    
	    instructions[20] = 32'b10001100000000010000001111101100;// lw r1,r0,1004
	    instructions[21] = 32'b00000000011000010001000000101010;// slt r2,r3,r1
	    instructions[22] = 32'b00000000000000000000000000000000;// nop
	    instructions[23] = 32'b00010000000000100000000000000001;// beq r2,r0,1
	    instructions[24] = 32'b00000000000000010001100000100000;// add r3,r1,r0
	    
	    instructions[25] = 32'b10001100000000010000001111101101;// lw r1,r0,1005
	    instructions[26] = 32'b00000000011000010001000000101010;// slt r2,r3,r1
	    instructions[27] = 32'b00000000000000000000000000000000;// nop
	    instructions[28] = 32'b00010000000000100000000000000001;// beq r2,r0,1
	    instructions[29] = 32'b00000000000000010001100000100000;// add r3,r1,r0
	    
	    instructions[30] = 32'b10001100000000010000001111101110;// lw r1,r0,1006
	    instructions[31] = 32'b00000000011000010001000000101010;// slt r2,r3,r1
	    instructions[32] = 32'b00000000000000000000000000000000;// nop
	    instructions[33] = 32'b00010000000000100000000000000001;// beq r2,r0,1
	    instructions[34] = 32'b00000000000000010001100000100000;// add r3,r1,r0
	    
	    instructions[35] = 32'b10001100000000010000001111101111;// lw r1,r0,1007
	    instructions[36] = 32'b00000000011000010001000000101010;// slt r2,r3,r1
	    instructions[37] = 32'b00000000000000000000000000000000;// nop
	    instructions[38] = 32'b00010000000000100000000000000001;// beq r2,r0,1
	    instructions[39] = 32'b00000000000000010001100000100000;// add r3,r1,r0
	    
	    instructions[40] = 32'b10001100000000010000001111110000;// lw r1,r0,1008
	    instructions[41] = 32'b00000000011000010001000000101010;// slt r2,r3,r1
	    instructions[42] = 32'b00000000000000000000000000000000;// nop
	    instructions[43] = 32'b00010000000000100000000000000001;// beq r2,r0,1
	    instructions[44] = 32'b00000000000000010001100000100000;// add r3,r1,r0
	    
	    instructions[45] = 32'b10001100000000010000001111110001;// lw r1,r0,1009
	    instructions[46] = 32'b00000000011000010001000000101010;// slt r2,r3,r1
	    instructions[47] = 32'b00000000000000000000000000000000;// nop
	    instructions[48] = 32'b00010000000000100000000000000001;// beq r2,r0,1
	    instructions[49] = 32'b00000000000000010001100000100000;// add r3,r1,r0
	    
  end
  assign instruction = instructions[address[15:2]];
endmodule

