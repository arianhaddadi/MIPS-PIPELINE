module Pipeline(input clk, rst);
	
	wire ID_PCLD, ID_IFTOIDREGLOAD, MEM_REGWRITE, EX_MEMREAD,EX_MEMREAD_OUT, ID_REGWRITE, ID_MEMREAD, ID_MEMWRITE, 
		 ID_MEMTOREG, ID_REGDST, ID_ALUSRC, ID_FLUSH, EX_REGWRITE, EX_MEMWRITE,EX_MEMWRITE_OUT, EX_MEMTOREG,EX_MEMTOREG_OUT,
		 EX_REGDST, EX_ALUSRC, EX_REGWRITE_OUT, WB_REGWRITE_OUT,WB_REGWRITE, MEM_REGWRITE_OUT,MEM_MEMREAD, MEM_MEMWRTIE,MEM_MEMTORREG,
		 MEM_MEMTORREG_OUT,WB_MEM_TO_REG   ;


	wire [1:0] ID_PCSRC;
	wire [4:0] MEM_RD, EX_RT,EX_RT_OUT, ID_RS, ID_RT, ID_RD, EX_RD, EX_RD_OUT, EX_RS, MEM_DEST_OUT,MEM_RD_OUT,WB_DEST_OUT, EX_DEST, MEM_DEST,WB_DEST;
	wire [5:0] ID_OPCODE, ID_FUNC,EX_FUNC, EX_OPCODE;
	wire [31:0] ID_JADDRESS, ID_BRANCH_ADDRESS, ID_PC_ADDED, IF_PC_ADDED, IF_INSTRUCTION, ID_INSTRUCTION,
				WB_WRITEDATA, MEM_ADDRESSORRES_OUT, MEM_ADDRESSORRES, ID_DATAREAD1, ID_DATAREAD2, ID_EXTENDED,EX_DATAREAD1, 
				EX_DATAREAD2,EX_EXTENDED, EX_RES, EX_B, MEM_DATA, MEM_MEMOUT, WB_RES, WB_DATA;

	IF instf(clk, rst, ID_PCLD, ID_PCSRC,ID_JADDRESS, ID_BRANCH_ADDRESS,/*Separator*/ IF_PC_ADDED, IF_INSTRUCTION);

	IFtoIDReg iftoidreg(clk, rst, ID_FLUSH, ID_IFTOIDREGLOAD, IF_INSTRUCTION, IF_PC_ADDED,/*Separator*/ ID_INSTRUCTION, ID_PC_ADDED);

	ID id(clk, rst, WB_REGWRITE, EX_MEMREAD_OUT,
	   	  MEM_RD_OUT, WB_DEST_OUT, EX_RT_OUT, 
	   	  MEM_ADDRESSORRES_OUT, ID_INSTRUCTION, ID_PC_ADDED, WB_WRITEDATA, /*Separator*/ 
	   	  ID_PCLD, ID_REGWRITE, ID_MEMREAD, ID_MEMWRITE, ID_MEMTOREG, ID_REGDST, ID_ALUSRC, ID_FLUSH, ID_IFTOIDREGLOAD,
	   	  ID_PCSRC,
	   	  ID_RS, ID_RD, ID_RT, 
	   	  ID_OPCODE, ID_FUNC,
	   	  ID_DATAREAD1, ID_DATAREAD2, ID_EXTENDED, ID_BRANCH_ADDRESS, ID_JADDRESS);	
		
	IDtoEXReg idtoexreg(clk, rst, ID_REGWRITE, ID_MEMREAD, ID_MEMWRITE, ID_MEMTOREG, ID_REGDST, ID_ALUSRC,
			  ID_DATAREAD1, ID_DATAREAD2, ID_EXTENDED,
			  ID_FUNC, ID_OPCODE,
			  ID_RS, ID_RT, ID_RD,/*Separator*/
			  EX_REGWRITE, EX_MEMREAD,  EX_MEMWRITE, EX_MEMTOREG, EX_REGDST, EX_ALUSRC,
			  EX_DATAREAD1, EX_DATAREAD2,EX_EXTENDED,
			  EX_FUNC, EX_OPCODE,
			  EX_RS, EX_RT, EX_RD);

	EX ex(EX_MEMREAD, EX_MEMWRITE, EX_REGWRITE, WB_REGWRITE_OUT, MEM_REGWRITE_OUT, EX_MEMTOREG, EX_REGDST, EX_ALUSRC,
	   EX_RD, EX_RS, EX_RT, MEM_DEST_OUT, WB_DEST_OUT,
	   EX_FUNC, EX_OPCODE,
	   EX_DATAREAD1, EX_DATAREAD2, EX_EXTENDED, MEM_ADDRESSORRES_OUT, WB_WRITEDATA,/*Separator*/
	   EX_MEMREAD_OUT, EX_MEMWRITE_OUT, EX_MEMTOREG_OUT, EX_REGWRITE_OUT, 
	   EX_RD_OUT, EX_DEST, EX_RT_OUT, 
	   EX_RES, EX_B);

	EXtoMEMReg extomemreg(clk, rst, EX_REGWRITE_OUT, EX_MEMREAD_OUT, EX_MEMWRITE_OUT, EX_MEMTOREG_OUT,
			   EX_RES, EX_B,
			   EX_RD_OUT, EX_DEST,/*Separator*/
			   MEM_REGWRITE, MEM_MEMREAD, MEM_MEMWRTIE, MEM_MEMTORREG,
			   MEM_ADDRESSORRES, MEM_DATA,
			   MEM_RD, MEM_DEST);

	MEM mem(clk, MEM_REGWRITE, MEM_MEMTORREG, MEM_MEMREAD, MEM_MEMWRTIE,
		MEM_RD, MEM_DEST,
		MEM_ADDRESSORRES, MEM_DATA,/*Separator*/
		MEM_REGWRITE_OUT, MEM_MEMTORREG_OUT, 
		MEM_DEST_OUT, MEM_RD_OUT,
		MEM_MEMOUT, MEM_ADDRESSORRES_OUT);

	MEMtoWBReg memtowbreg(clk, rst, MEM_REGWRITE_OUT, MEM_MEMTORREG_OUT,
				MEM_ADDRESSORRES_OUT, MEM_MEMOUT,
				MEM_DEST_OUT,/*Separator*/
				WB_REGWRITE, WB_MEM_TO_REG,
				WB_RES, WB_DATA,
				WB_DEST);

	WB wb(WB_REGWRITE, WB_MEM_TO_REG, WB_DEST,WB_DATA, WB_RES, /*Separator*/WB_REGWRITE_OUT, WB_DEST_OUT, WB_WRITEDATA);

endmodule



